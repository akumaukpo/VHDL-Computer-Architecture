library ieee;
use ieee.std_logic_1164.all;

package special is
  type twod_arr is array ( integer range<> , integer range<> ) of std_logic;
end special;
